
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY rom_block IS
   PORT (addra: IN std_logic_VECTOR(9 DOWNTO 0);
         addrb: IN std_logic_VECTOR(9 DOWNTO 0);
         clka:  IN std_logic;
         clkb:  IN std_logic;
         douta: OUT std_logic_VECTOR(15 DOWNTO 0);
         doutb: OUT std_logic_VECTOR(15 DOWNTO 0);
         ena:   IN std_logic;
         enb:   IN std_logic);
END rom_block;

library unisim;
use unisim.vcomponents.all;

architecture low_level_definition of rom_block is

begin

-- The synchronous set/reset input, SSR, forces the data output latches to value specified by the
-- SRVAL attribute. When SSR and the enable signal, EN, are High, the data output latches for
-- the DO and DOP outputs are synchronously set to a '0' or '1' according to the SRVAL parameter.

   --Instantiate the Xilinx primitive for a block RAM
   u1: RAMB16_S18_S18
   --INIT values repeated to define contents for functional simulation
   generic map( INIT_A  => X"00000",
                INIT_B  => X"00000",
                SRVAL_A => X"00000",
                SRVAL_B => X"00000",
                INIT_00 => X"FFD2FFC8FFDB001100130044003CFFA1FFB9000CFFA90021003800190063FFD7",
                INIT_01 => X"003F0052FFBBFFB8FFE700400048000A001BFFE5FFAFFFB6004600260013FFC8",
                INIT_02 => X"0028FFE6001D0047FFD90060FFEB0011FFB9FFF1000A0010FFB2FFBB0016FFCB",
                INIT_03 => X"0061002CFFC9FFE90023000EFFF1FFEB001BFFD9FFB2FFF5FFF40056FFF3FFF2",
                INIT_04 => X"0062005D004B000AFFC6000BFFE2001E0045FFCC0061001000180012004CFFE5",
                INIT_05 => X"FFA3FFB0FFDAFFEF0014FFBA0025FFE6FFD3FFA7FFC9000EFFD90026FFA70012",
                INIT_06 => X"FFCD005D00300055000B003CFFE0FFE80040FFC00027FFD30062FFCAFFDFFFE4",
                INIT_07 => X"003DFF9DFFAF004EFFC40021FFA50017FFCA004FFFB3FFEBFFB50037001A001A",
                INIT_08 => X"FFA7FFA6004E00130016FFA40013FFF0FFDDFFF10063000F002CFFA30021FFF4",
                INIT_09 => X"FFC9FFB3002EFFDA000D00380030003E0048FFB10030002300490049FFA80024",
                INIT_0A => X"000BFFEFFFCFFFDD0056005DFFE5FFB90054FFF30011FFB10036005EFFA5FFF6",
                INIT_0B => X"FFA2FFB2FFA10054FFB2000FFFEA00190035FFF0001EFFD70054001C0011FFED",
                INIT_0C => X"FFC100150010FFF6FFDE0027005900170061FFB3FFF3004C0032FFBAFFE4FFC1",
                INIT_0D => X"FFE0005B003F0017FFDEFFE0002B00100051FFA0FFE3FFC8FFC8000D0015FFF2",
                INIT_0E => X"0027FFBAFFC0FFF5000FFFC2FFDEFFCAFFE1FFF0FFC80022FF9E0013FF9EFFD5",
                INIT_0F => X"FFB80012FFA1000F000BFFABFFBCFFF0FFA3FFAEFFF4FFB7FFCF002E00110021",
                INIT_10 => X"0016FFED0050001000260056005CFFE6FFD5FFE40063001B00120052FFC7001B",
                INIT_11 => X"0042FFA80056FFE7FFE1FFF1FFE90024FFEBFFAC005DFF9DFF9FFFF40015FFAE",
                INIT_12 => X"004AFFEE0014003CFFF3FFB8005B0029FFBF00590046FFF1FFD2000A0046004B",
                INIT_13 => X"0039FFED000C0010FFAF0044000BFFBF001BFFC20012004C0038FFE4003E000B",
                INIT_14 => X"FFE5001B0012000D0038002D0050004AFFF5FFC90045FFA9FFF1002F004FFFC5",
                INIT_15 => X"0027001C00120019FFEF000A001D0020FFCEFFBB000B002AFFE0FFF5001DFFD2",
                INIT_16 => X"FFD70031FFEC000CFFE1000FFFDA0056000C000D0020001AFFC8000B00340035",
                INIT_17 => X"FFCEFFF0FFBD003CFFB1000B000C00110024000AFFDDFFF500110054FFA1002E",
                INIT_18 => X"FFE2000E0047000A004A004C001500480011000FFFDEFFF4FFF3000E0024005C",
                INIT_19 => X"FFEDFFCE0038FFBF001FFFEBFFC8003400430033FFAA000B005DFFD00048004F",
                INIT_1A => X"FFC5001CFFF6FFB000330013000B001FFFD200110012000AFFB700320048FFE5",
                INIT_1B => X"FFBC0012001FFFE10034FFEC005D000DFFEAFFF6003400570010FFCDFFD4000B",
                INIT_1C => X"0040000E0037000F005DFFB5FFABFFDFFFED004EFFA4000D000AFFC7FFECFFCC",
                INIT_1D => X"FFEDFFA8003200610016FFDCFFA50061FFDA0014FFC5FFF5FFE8000D00190025",
                INIT_1E => X"0014004F000E00200015FFC4FFA40018FFEDFFE1002800520012FFE2FFEEFFB3",
                INIT_1F => X"000B0025FFCE005BFFC80029000AFFE1002FFFB40019000E0034004F005DFFEC",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_00 => X"3CCCCFC0C00F333FFF33FCCC00CC30030F0F3FCF30CCF0F30FC03F03FC03CC03",
               INITP_01 => X"FCCC33033F0F330FF300300CF033F0333CCCCFC0C00F333FFF33FCCC00CC3003",
               INITP_02 => X"CC3FFFC03F3FFCCFC0F03FC3C3C03C3FFCCC33033F0F330FF300300CF033F033",
               INITP_03 => X"30C3303030F0C3C033FCF3F33003F00CCC3FFFC03F3FFCCFC0F03FC3C3C03C3F",
               INITP_04 => X"FCC00F0CCCCC00C000C0F0F3C000F3C330C3303030F0C3C033FCF3F33003F00C",
               INITP_05 => X"C330F03CCF00C0C3F33C0C30C0000FC0FCC00F0CCCCC00C000C0F0F3C000F3C3",
               INITP_06 => X"0CC33003003CF03FF03CCFC0003FCC3FC330F03CCF00C0C3F33C0C30C0000FC0",
               INITP_07 => X"000000000000000000000000000000000CC33003003CF03FF03CCFC0003FCC3F")

     PORT MAP (DOA   => douta,
               DOB   => doutb,
               DOPA  => open,
               DOPB  => open,
               ADDRA => addra,
               ADDRB => addrb,
               CLKA  => clka,
               CLKB  => clkb,
               DIA   => (OTHERS => '0'),
               DIB   => (OTHERS => '0'),
               DIPA  => (OTHERS => '0'),
               DIPB  => (OTHERS => '0'),
               ENA   => ena,
               ENB   => enb,
               SSRA  => '0',
               SSRB  => '0',
               WEA   => '0',
               WEB   => '0');


end low_level_definition;

